`define INSTR_MEM_FILE "tests/b_instr.mem"
`define DATA_MEM_FILE "tests/b_data.mem"
`define MAX_CYCLES 2000
