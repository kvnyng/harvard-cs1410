`define INSTR_MEM_FILE "tests/rtype_tests_instr.mem"
`define DATA_MEM_FILE ""
`define MAX_CYCLES 2000
