`define INSTR_MEM_FILE "tests/c_instr.mem"
`define DATA_MEM_FILE "tests/c_data.mem"
`define MAX_CYCLES 2000
