module and32
    (
        input logic [31:0] x, [31:0] y,
        output logic [31:0] z
    );

    // TODO: Implement the AND gate output. 
    //       Hint: the code is very short, this is 
    //       just to show you how module heirarchy works. 

    // YOUR CODE HERE
    assign z = 0;

endmodule
