`timescale 1ns / 1ps

module timer
    #(parameter N = 5)
    (
        input logic clk, clk_slow,
        input logic rst, en, load,
        input logic [N-1:0] init,
        output logic [N-1:0] out
    );

    /*** IMPORTANT NOTE ********************************************************
    * Please make sure to write your synchronous always blocks as such:

    always_ff @(posedge clk, posedge rst) begin
        if (rst) begin
            // asynchronous reset
        end
        else if (clk_en) begin
            // do stuff
        end
    end

    * or as such:

    always_ff @(posedge clk) begin
        if (rst) begin
            // synchronous reset
        end
        else if (clk_en) begin
            // do stuff
        end
    end

    * where clk is the 100 MHz system clock and clk_en is the 1 Hz "clock"
    * produced by your clock divider.
    *
    * Why is this the correct way to write things? Behind the scenes, clk is
    * generated by specialized clock generation circuitry within the FPGA chip,
    * while clk_en (the 1 Hz "clock") is not. This means that clk_en will be a
    * VERY bad choice of signal to clock FFs with and may cause a slew of subtle
    * bugs -- it's not a "real" clock. Additionally, directly clocking FFs with
    * such slow clocks is NEVER a good idea for lots of lower level electronics
    * reasons.
    *
    * If you put the 1 Hz "clock" in the sensitivity list of an always block,
    * you will lose points. So don't do it.
    *
    * Bug Jon if you're curious and want to know more.
    ***************************************************************************/

    // implements the timer specified in the lab guide
    
     always_ff @(posedge clk) begin
        if (rst) begin
            out <= 5'd0;  // Start at 0, not 15
        end
        else if (load) begin
            out <= init;  // Load the initial value
        end
        else if (en & clk_slow & out != 0) begin
            out <= out - 1;        
        end
    end

endmodule
