module cla
    (
         // inputs/outputs here
    );

    // TODO (part 2): implement carry-lookahead adder
    //       Be sure to comment out the module instantiation 
    //       of your old ripple-carry adder in STUDENT_alu.sv

endmodule
