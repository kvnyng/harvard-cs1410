// SV Header for ALU op-codes
// Use in your code with: `opcode, for example `ALU_ADD
`define ALU_AND 3'b000
`define ALU_ADD 3'b001
`define ALU_SUB 3'b010
`define ALU_SLT 3'b011
`define ALU_SRL 3'b100
`define ALU_SRA 3'b101
`define ALU_SLL 3'b110
