module sra
    (
         // inputs/outputs here
    );

    // TODO (part 2): implement sra

endmodule
