module slt
    (
         // inputs/outputs here
    );

    // TODO: implement slt

endmodule
