module adder
    (
         // inputs/outputs here
    );

    // TODO: implement adder

endmodule
