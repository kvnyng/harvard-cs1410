module sll
    (
         // inputs/outputs here
    );

    // TODO (part 2): implement sll

endmodule
