module srl
    (
         // inputs/outputs here
    );

    // TODO (part 2): implement srl

endmodule
